PK   P�S��g)      cirkitFile.json�]]o����+�^�W���$y�N��h��)rs`�D5B}$W��A�{�Kږ�_�<'r.��yv�zv8;�~X������xn�N��a�Nȫշ�i�}y��Z�������O����w?������C�9~�?���ֈ��^Wk�L���T���ծ�P}�6��z�����OV������1u��[L���[L�i��� �'@�	�z� �'@�	�~��'Q���Ӯe�z��Tj+6�ZF��l7�6��g#C+dh	�C�AY��j�èmk�F�նn��n�M���Udh�mb�6C�m%��띭�����f�m6�z�=x�24v��
��
W�
W��*�ئ7� �y����e��]���Mo�*W����ӷ7�z��FRO��H��{I=}k#���l$�4�I�i��h���]&������U4}�{�����/W��A�e�*�>��@�I��_2LѶ_�۝�d3�ڲ_W�M�T��Z�c�����6t*L!-��Sa
i�T�D\0>L�F�ͺ�vRW���h��U�֢��]�כ]�h��p~��
Z CC4Uhh���PL�h�R۟��۝���Z�Jo�Puf�T}#����`۝c*2vʱ��� ��
[$�il��n���e��K��!�� @�A�]�F�?`�� T�A��P�S5����g@�t��π�3 ��?�ς�� �,�?���|�z��i�
�^{z���+���^x$���#���I=��h�Ai�.�����ˤ�h� �2�/�>ȾLꋦ�/����~�_&�E��'A�I��L����d��n��@n��457����CQs�ةG��� 2v*�E� c��\��\��\��\���g2��>x��dWh�h��/�]����dWh� �2���_&�B���ɮ���-ȿLv���/�]����dWh� �2��~��g���?� ����:R�����S�q�OJ��SO�HC�]I=�iH�iGCRO��K��i��_���wd˓˄2tڷ_�E,OmaIC����.byjL:O�^�E,On�)Cg��˓�o���9'�2��CS�_�B�N}���Ð��5�ە�m�w�Xv�����[E��Z}ƀ"YP�fA1,(��aAiYP:�1�������������������Â�Ă�Œ�Œ�{�v(�g�}�J�%�y��,6���F`,�5��>4��B`xX,yX�xX��,�}1���R�-P+�P�7j]J�@�c@).%j������rTC�'��!p9�!�q��p�Ր+�8���Q����Œ��ST�S[3��,��r��x�1����x�jr����Y#����"�N5���\r�J�XcsrA�gqg�Z�G`f_l>��i�/�kSK��k_�y|��a�f��y|��(4OD�y"
��5������Ǝ�ņ�ņ�ņ�ņ�Ŗ�Ŗ�Ŗ�Ŷ�bj�Jqf��K(<�R\�Ԓ&��Ҧ81�6�܉�uL��ao9kC.���!p9kC�����p9kC.���z<,.gmȕT0<,.gm��U0<,�<,��6�M<�|�f���r䢦|.�\����K�8"++++_\�ڐ�8`x|q9kC.:��aq9kC�D��aq9kC.O��u𰸜�!�,q�𰸜�!2q�𰸜�!W7q�𰸜�!�<q�𰸜���A�c6jI�-����Zh��G�b���ڦV1�W6����bi�-�/����>y[�5?�y���0���%��$� �ঈu9�=!�Ć��ٿ��ܤ��m����߷����_��V�<���R��p��Z�rϧ�.n�8G�,(�E��˂Ұ��,(����^�C_��_�C`��`�Ca��a�Cb��b��b��yX,yX,yX,yX,yX,yX,yX,yX�xX��,&��(<��8G).'rq
�R\L�������)�c"/{�Q�8����娆^�� ���rTC/Na�z<,.G5����zq
��Q�8����娆^�� �J�X�X�X�X�X�X�X�X�X�X3E�<,�<,�<,�<,�<,�<,6<,6<,6<,6<,6L;[[[�"���)8Jqf��)8
ϼ7�8G).mrq
�R\����1������8������8������8���񰸜���0�𰸜���0�𰸜���0�𰸜���0�0�<,.gm��)0<,.gm��)0<,.gm��)0<,.gm��)0<,.gm��)0<,.gm��)0<,.gm��)0L;��6����6����6��,�8G)��8Gᙗ��&��(ťM.NɣP�Sp�2_��)8J�/���8/���|����(e�K-N�Q��B.N�Q��B.NyB��j��_��wSn����Iq��~n���Ͱ��n���pZ����0�����~GJs@cC�26v���	��n�d4v��/5���@o!C'J��N!C�'dh�+rbhj��@C'xFꠡ��7AC'91L�_���'�ł�Щ-�KM� �b��G���9�fus�6�����Ƹ�?lc!���_0��q�c&��$�	hT�`\2��Ƙ&��fք7�8q��� �?q�04k��D��A)�`��`'z�����mz� �ȿ��d�/�-��3��, C��o���=n׻Ⱦ?m���Fϟ�����=�hw�[�{P_��
�נ��-�߀�-�ߡ��	�2P�(JB��P�4(JD�2Q�L��/tL�_��[����<�ǣM���6�KD��6D�D�K�G�B9�2'�B���3Ξ�e�ϸzrg!D?���݄�� w��e`.ޠw
� P��z_  �a.ޠw�<��\�A���L�(c!�;��DB���g��254a]`P��p�!���*���5��0���z=�	W@�z���x�Ϙ�!�,,� ��FݺFݺF)�� u�04`h4�Ш��h�aP&��e�A�h���D�2ѠL4(�D�2ѢL�(m����=�~f��z}��3�ܜ��,CrCD?��Mx ��D�K|Л�@ (	s�zk �a.�Ao�y"�����m�21���7Ɂ P&J��2�������7ɡ���rh;az��N��?���7ҁB��
�B9�Po�Po��G���@ ����#��p  ���|���21���7�� P&����6 �B���G���@ (s�z� eb.AoM�  7�Y��ρ��ip��$�65��S r��\�!�q2��5LnV��gV0�A�"�N��N5�9����cά,r���9���ܯ1'2;���ܲ&帨�j�6AԮ5�9��I��k�[�,�AXy��{�&68�S�/0���I�\Q��ջO+�Z�q�tK��}��;{����_���x
�e���3�⇿>?g�iH�!=����z�J�+�j_0#��t�i�� +ʃ�_����9N×o�j_9�+x}%��h�NC;�4������v�ih����q�i�a����4��0N�8�4�ӰN�:뺏�(q�o�����	���n�!ШH��D)�6�H�b�oF��8y��pvN�v<�]��S���Ҥ�92n��	s�n]a1n�&ys��^a1n�����M�p[X7�Ѐ5p�0? X��xqkަ�X��E�A��<���V��E�Aq��M��7W��D�A�u����5o��+ܪ��M��}8`��%J=�αw�z�s���C������n��D�"��,��H�"��,ҡ��"��,����EM(jgQ��Y�"�4"��<�|���ᄈ�	ገ�ᔈ�)ᜈ�9ᤈ�Iᬈ�Y�����ݮOC�]�����;���Ύ���������9��mF�0rt�UJ�v��f{kG�����8��F]������ߜ�Ǹ�H=|՟��诧��p:���|p�sa4��|��>^ڡ��>;������}���o*1�ss�x؏ìƿ�=~��×#��ݮ�{F��p�f��_���N�?��a�zw�i�����q�oΏ'�/m��i/�|��O���x`0e�����?��T|�B^�+U�q�Iغ,�#'�몺^7U�i�U?F��V5V�M۹��?<���f�!eۮV��~���i���Vǯn�����I�Ѥ�o_]I�\�FE�L����I-%�ZzҒ����H6�xȩ�]Z����j'0�K���hS]B��Q��৿�>�m^#�����9틮���oe^Ι�n.���q}q���/`D.y��4�i��1¯�	n<y��?<?n��o����lq]_ףcD�P�]�/�~�o���q�����/��UR����++�_8/��*�ݍ��m���YwM�v��Z��n�`v��,=)���L���_���2�[ʕ��Z��vH�][UkafA3J��,��5���Z�X�ʄ�i�n�hl*�P�`���1�է���a:M�����t��a>M]��.OS����A��i�rPk_J(��C��^��^��^������&!P)�Ҩ����j�U�Ni���Hi�	�٪.eUDФ4�i�+o�VL2��$3�\���-�$3ZD2��ŷ��b�-"�њ$ZD2�E$3ZkShɌ�̮�N���N""��Dʶ�dF�HF��nÌ���]�a���nâ"��λ�m3�u}�lgZ�r��rd����d�"m��xxZ���Q	��`��&(��*"��"�	J���&��`�j�e�P�x�.q}��(r��S�9�q"�=�m�8��'r���uE��[s�J�/����۲Z\p�lOp\'�W��E��:~�l�I�o�O��g�����pd����p�=��	'<�qd��"g��q�9>��'<>��'� tL0!E�J8��`�������_E�M����W�7��'�^ �փ�æ2��ԪR��Ͷ���W[��� ��Je��K
i]�=��4�T{!Qͥ�4����%�>!�I���i�׿}��|���+�ş>|�P�����/�S��l4�#c�1�+��릩��Kb���U��m�m5��1����c�j�ݺ�Ȕ�)u�[��lI̔��O��Z_F>���P��ނJZu�J�K�E�Dz�𿠒��f���~��/�2ыR ��Yo¬V�bV�2��V�ì��IM�ǻ.E�@�S�����J����/?�#��(9z��H��Mu���Z�FwV���Z�dյͶR�0T�ںi����CY�ɤ�KOW��I��)Ic�����?PK
   P�S��g)                    cirkitFile.jsonPK      =   V    